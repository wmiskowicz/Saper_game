`timescale 1ns / 1ps
// ROM with synchonous read (inferring Block RAM)
// character ROM
//  - 8-by-16 (8-by-2^4) font
//  - 128 (2^7) characters
//  - ROM size: 512-by-8 (2^11-by-8) bits
//              16K bits: 1 BRAM

module num_font_rom
    (
        input  wire        clk,
        input  wire [11:0] addr,            // {char_code[5:0], char_line[5:0]}
        output reg  [49:0]  char_line_pixels, // pixels of the character line
        output reg  [11:0] num_color
    );
    import colour_pkg::*;

    // body
    always_ff@(posedge clk)begin
        case(addr[11:6])
            6'h31: num_color <= NUM_1;
            6'h32: num_color <= NUM_2;
            6'h33: num_color <= NUM_3;
            6'h34: num_color <= NUM_4;
            6'h35: num_color <= NUM_5;
            6'h36: num_color <= NUM_6;
            6'h37: num_color <= NUM_7;
            default: num_color <= NUM_DEFAULT;
        endcase

        case (addr)
            //code x00
            12'h000: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h001: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h002: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h003: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h004: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h005: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h006: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h007: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h008: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h009: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h00a: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h00b: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h00c: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h00d: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h00e: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h00f: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h010: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h011: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h012: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h013: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h014: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h015: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h016: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h017: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h018: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h019: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h01a: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h01b: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h01c: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h01d: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h01e: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h01f: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h020: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h021: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h022: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h023: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h024: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h025: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h026: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h027: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h028: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h029: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h02a: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h02b: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h02c: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h02d: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h02e: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h02f: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h030: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'h031: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            
            
            //code x31
            12'hc40: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc41: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc42: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc43: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc44: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc45: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc46: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc47: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc48: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc49: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc4a: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc4b: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc4c: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc4d: char_line_pixels <= 50'b00000000000000000000000111100000000000000000000000; //
            12'hc4e: char_line_pixels <= 50'b00000000000000000000000111100000000000000000000000; //
            12'hc4f: char_line_pixels <= 50'b00000000000000000000011111100000000000000000000000; //
            12'hc50: char_line_pixels <= 50'b00000000000000000000011111100000000000000000000000; //
            12'hc51: char_line_pixels <= 50'b00000000000000000001111111100000000000000000000000; //
            12'hc52: char_line_pixels <= 50'b00000000000000000001111111100000000000000000000000; //
            12'hc53: char_line_pixels <= 50'b00000000000000000000000111100000000000000000000000; //
            12'hc54: char_line_pixels <= 50'b00000000000000000000000111100000000000000000000000; //
            12'hc55: char_line_pixels <= 50'b00000000000000000000000111100000000000000000000000; //
            12'hc56: char_line_pixels <= 50'b00000000000000000000000111100000000000000000000000; //
            12'hc57: char_line_pixels <= 50'b00000000000000000000000111100000000000000000000000; //
            12'hc58: char_line_pixels <= 50'b00000000000000000000000111100000000000000000000000; //
            12'hc59: char_line_pixels <= 50'b00000000000000000000000111100000000000000000000000; //
            12'hc5a: char_line_pixels <= 50'b00000000000000000000000111100000000000000000000000; //
            12'hc5b: char_line_pixels <= 50'b00000000000000000000000111100000000000000000000000; //
            12'hc5c: char_line_pixels <= 50'b00000000000000000000000111100000000000000000000000; //
            12'hc5d: char_line_pixels <= 50'b00000000000000000000000111100000000000000000000000; //
            12'hc5e: char_line_pixels <= 50'b00000000000000000000000111100000000000000000000000; //
            12'hc5f: char_line_pixels <= 50'b00000000000000000000111111111100000000000000000000; //
            12'hc60: char_line_pixels <= 50'b00000000000000000001111111111110000000000000000000; //
            12'hc61: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc62: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc63: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; // 
            12'hc64: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc65: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc66: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc67: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc68: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc69: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc6a: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc6b: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc6c: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc6d: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc6e: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc6f: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc70: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc71: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //


            //code x32
            12'hc80: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc81: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc82: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc83: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc84: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc85: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc86: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc87: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc88: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc89: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc8a: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc8b: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc8c: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hc8d: char_line_pixels <= 50'b00000000000000000001111111111000000000000000000000; //
            12'hc8e: char_line_pixels <= 50'b00000000000000000011111111111100000000000000000000; //
            12'hc8f: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'hc90: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'hc91: char_line_pixels <= 50'b00000000000000000000000000011110000000000000000000; //
            12'hc92: char_line_pixels <= 50'b00000000000000000000000000111100000000000000000000; //
            12'hc93: char_line_pixels <= 50'b00000000000000000000000001111000000000000000000000; //
            12'hc94: char_line_pixels <= 50'b00000000000000000000000011110000000000000000000000; //
            12'hc95: char_line_pixels <= 50'b00000000000000000000000111100000000000000000000000; //
            12'hc96: char_line_pixels <= 50'b00000000000000000000001111000000000000000000000000; //
            12'hc97: char_line_pixels <= 50'b00000000000000000000011110000000000000000000000000; //
            12'hc98: char_line_pixels <= 50'b00000000000000000000111100000000000000000000000000; //
            12'hc99: char_line_pixels <= 50'b00000000000000000001111000000000000000000000000000; //
            12'hc9a: char_line_pixels <= 50'b00000000000000000011110000000000000000000000000000; //
            12'hc9b: char_line_pixels <= 50'b00000000000000000111100000000000000000000000000000; //
            12'hc9c: char_line_pixels <= 50'b00000000000000000111100000000000000000000000000000; //
            12'hc9d: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'hc9e: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'hc9f: char_line_pixels <= 50'b00000000000000000111111111111110000000000000000000; //
            12'hca0: char_line_pixels <= 50'b00000000000000000111111111111110000000000000000000; //
            12'hca1: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hca2: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hca3: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; // 
            12'hca4: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hca5: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hca6: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hca7: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hca8: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hca9: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hcaa: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hcab: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hcac: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hcad: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hcae: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hcaf: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hcb0: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hcb1: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //


            //code x33
            12'hcc0: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hcc1: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hcc2: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hcc3: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hcc4: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hcc5: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hcc6: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hcc7: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hcc8: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hcc9: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hcca: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hccb: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hccc: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hccd: char_line_pixels <= 50'b00000000000000000001111111111000000000000000000000; //
            12'hcce: char_line_pixels <= 50'b00000000000000000011111111111100000000000000000000; //
            12'hccf: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'hcd0: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'hcd1: char_line_pixels <= 50'b00000000000000000000000000011110000000000000000000; //
            12'hcd2: char_line_pixels <= 50'b00000000000000000000000000011110000000000000000000; //
            12'hcd3: char_line_pixels <= 50'b00000000000000000000000000011110000000000000000000; //
            12'hcd4: char_line_pixels <= 50'b00000000000000000000000000111100000000000000000000; //
            12'hcd5: char_line_pixels <= 50'b00000000000000000000011111111000000000000000000000; //
            12'hcd6: char_line_pixels <= 50'b00000000000000000000011111111000000000000000000000; //
            12'hcd7: char_line_pixels <= 50'b00000000000000000000000000111100000000000000000000; //
            12'hcd8: char_line_pixels <= 50'b00000000000000000000000000011110000000000000000000; //
            12'hcd9: char_line_pixels <= 50'b00000000000000000000000000011110000000000000000000; //
            12'hcda: char_line_pixels <= 50'b00000000000000000000000000011110000000000000000000; //
            12'hcdb: char_line_pixels <= 50'b00000000000000000000000000011110000000000000000000; //
            12'hcdc: char_line_pixels <= 50'b00000000000000000000000000011110000000000000000000; //
            12'hcdd: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'hcde: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'hcdf: char_line_pixels <= 50'b00000000000000000011111111111100000000000000000000; //
            12'hce0: char_line_pixels <= 50'b00000000000000000001111111111000000000000000000000; //
            12'hce1: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hce2: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hce3: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; // 
            12'hce4: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hce5: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hce6: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hce7: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hce8: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hce9: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hcea: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hceb: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hcec: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hced: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hcee: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hcef: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hcf0: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hcf1: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //


            //code x34
            12'hd00: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd01: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd02: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd03: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd04: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd05: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd06: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd07: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd08: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd09: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd0a: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd0b: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd0c: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd0d: char_line_pixels <= 50'b00000000000000000000000000111000000000000000000000; //
            12'hd0e: char_line_pixels <= 50'b00000000000000000000000001111000000000000000000000; //
            12'hd0f: char_line_pixels <= 50'b00000000000000000000000111111000000000000000000000; //
            12'hd10: char_line_pixels <= 50'b00000000000000000000000111111000000000000000000000; //
            12'hd11: char_line_pixels <= 50'b00000000000000000000011111111000000000000000000000; //
            12'hd12: char_line_pixels <= 50'b00000000000000000000011111111000000000000000000000; //
            12'hd13: char_line_pixels <= 50'b00000000000000000001111001111000000000000000000000; //
            12'hd14: char_line_pixels <= 50'b00000000000000000001111001111000000000000000000000; //
            12'hd15: char_line_pixels <= 50'b00000000000000000111100001111000000000000000000000; //
            12'hd16: char_line_pixels <= 50'b00000000000000000111100001111000000000000000000000; //
            12'hd17: char_line_pixels <= 50'b00000000000000000111111111111110000000000000000000; //
            12'hd18: char_line_pixels <= 50'b00000000000000000111111111111110000000000000000000; //
            12'hd19: char_line_pixels <= 50'b00000000000000000000000001111000000000000000000000; //
            12'hd1a: char_line_pixels <= 50'b00000000000000000000000001111000000000000000000000; //
            12'hd1b: char_line_pixels <= 50'b00000000000000000000000001111000000000000000000000; //
            12'hd1c: char_line_pixels <= 50'b00000000000000000000000001111000000000000000000000; //
            12'hd1d: char_line_pixels <= 50'b00000000000000000000000001111000000000000000000000; //
            12'hd1e: char_line_pixels <= 50'b00000000000000000000000001111000000000000000000000; //
            12'hd1f: char_line_pixels <= 50'b00000000000000000000000011111100000000000000000000; //
            12'hd20: char_line_pixels <= 50'b00000000000000000000000111111110000000000000000000; //
            12'hd21: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd22: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd23: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; // 
            12'hd24: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd25: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd26: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd27: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd28: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd29: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd2a: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd2b: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd2c: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd2d: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd2e: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd2f: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd30: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd31: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //


            //code x35
            12'hd40: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd41: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd42: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd43: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd44: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd45: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd46: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd47: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd48: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd49: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd4a: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd4b: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd4c: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd4d: char_line_pixels <= 50'b00000000000000000111111111111110000000000000000000; //
            12'hd4e: char_line_pixels <= 50'b00000000000000000111111111111110000000000000000000; //
            12'hd4f: char_line_pixels <= 50'b00000000000000000111100000000000000000000000000000; //
            12'hd50: char_line_pixels <= 50'b00000000000000000111100000000000000000000000000000; //
            12'hd51: char_line_pixels <= 50'b00000000000000000111100000000000000000000000000000; //
            12'hd52: char_line_pixels <= 50'b00000000000000000111100000000000000000000000000000; //
            12'hd53: char_line_pixels <= 50'b00000000000000000111100000000000000000000000000000; //
            12'hd54: char_line_pixels <= 50'b00000000000000000111100000000000000000000000000000; //
            12'hd55: char_line_pixels <= 50'b00000000000000000111111111110000000000000000000000; //
            12'hd56: char_line_pixels <= 50'b00000000000000000011111111111100000000000000000000; //
            12'hd57: char_line_pixels <= 50'b00000000000000000000000000011110000000000000000000; //
            12'hd58: char_line_pixels <= 50'b00000000000000000000000000011110000000000000000000; //
            12'hd59: char_line_pixels <= 50'b00000000000000000000000000011110000000000000000000; //
            12'hd5a: char_line_pixels <= 50'b00000000000000000000000000011110000000000000000000; //
            12'hd5b: char_line_pixels <= 50'b00000000000000000000000000011110000000000000000000; //
            12'hd5c: char_line_pixels <= 50'b00000000000000000000000000011110000000000000000000; //
            12'hd5d: char_line_pixels <= 50'b00000000000000000111000000011110000000000000000000; //
            12'hd5e: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'hd5f: char_line_pixels <= 50'b00000000000000000011111111111000000000000000000000; //
            12'hd60: char_line_pixels <= 50'b00000000000000000001111111110000000000000000000000; //
            12'hd61: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd62: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd63: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; // 
            12'hd64: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd65: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd66: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd67: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd68: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd69: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd6a: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd6b: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd6c: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd6d: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd6e: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd6f: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd70: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd71: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            

            //code x36
            12'hd80: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd81: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd82: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd83: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd84: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd85: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd86: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd87: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd88: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd89: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd8a: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd8b: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd8c: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hd8d: char_line_pixels <= 50'b00000000000000000000001111110000000000000000000000; //
            12'hd8e: char_line_pixels <= 50'b00000000000000000000111111100000000000000000000000; //
            12'hd8f: char_line_pixels <= 50'b00000000000000000001111100000000000000000000000000; //
            12'hd90: char_line_pixels <= 50'b00000000000000000011111000000000000000000000000000; //
            12'hd91: char_line_pixels <= 50'b00000000000000000111110000000000000000000000000000; //
            12'hd92: char_line_pixels <= 50'b00000000000000000111100000000000000000000000000000; //
            12'hd93: char_line_pixels <= 50'b00000000000000000111100000000000000000000000000000; //
            12'hd94: char_line_pixels <= 50'b00000000000000000111100000000000000000000000000000; //
            12'hd95: char_line_pixels <= 50'b00000000000000000111111111111000000000000000000000; //
            12'hd96: char_line_pixels <= 50'b00000000000000000111111111111100000000000000000000; //
            12'hd97: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'hd98: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'hd99: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'hd9a: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'hd9b: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'hd9c: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'hd9d: char_line_pixels <= 50'b00000000000000000111000000011110000000000000000000; //
            12'hd9e: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'hd9f: char_line_pixels <= 50'b00000000000000000011111111111100000000000000000000; //
            12'hda0: char_line_pixels <= 50'b00000000000000000001111111110000000000000000000000; //
            12'hda1: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hda2: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hda3: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; // 
            12'hda4: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hda5: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hda6: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hda7: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hda8: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hda9: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdaa: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdab: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdac: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdad: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdae: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdaf: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdb0: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdb1: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //


            //code x37
            12'hdc0: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdc1: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdc2: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdc3: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdc4: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdc5: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdc6: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdc7: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdc8: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdc9: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdca: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdcb: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdcc: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdcd: char_line_pixels <= 50'b00000000000000000111111111111110000000000000000000; //
            12'hdce: char_line_pixels <= 50'b00000000000000000111111111111110000000000000000000; //
            12'hdcf: char_line_pixels <= 50'b00000000000000000111110000111110000000000000000000; //
            12'hdd0: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'hdd1: char_line_pixels <= 50'b00000000000000000000000000011110000000000000000000; //
            12'hdd2: char_line_pixels <= 50'b00000000000000000000000000011110000000000000000000; //
            12'hdd3: char_line_pixels <= 50'b00000000000000000000000000011110000000000000000000; //
            12'hdd4: char_line_pixels <= 50'b00000000000000000000000000011110000000000000000000; //
            12'hdd5: char_line_pixels <= 50'b000000000000000000000000000111100000000000000000000; //
            12'hdd6: char_line_pixels <= 50'b00000000000000000000000001111000000000000000000000; //
            12'hdd7: char_line_pixels <= 50'b00000000000000000000000111100000000000000000000000; //
            12'hdd8: char_line_pixels <= 50'b00000000000000000000001111000000000000000000000000; //
            12'hdd9: char_line_pixels <= 50'b00000000000000000000011110000000000000000000000000; //
            12'hdda: char_line_pixels <= 50'b00000000000000000000011110000000000000000000000000; //
            12'hddb: char_line_pixels <= 50'b00000000000000000000011110000000000000000000000000; //
            12'hddc: char_line_pixels <= 50'b00000000000000000000011110000000000000000000000000; //
            12'hddd: char_line_pixels <= 50'b00000000000000000000011110000000000000000000000000; //
            12'hdde: char_line_pixels <= 50'b00000000000000000000011110000000000000000000000000; //
            12'hddf: char_line_pixels <= 50'b00000000000000000000011110000000000000000000000000; //
            12'hde0: char_line_pixels <= 50'b00000000000000000000011110000000000000000000000000; //
            12'hde1: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hde2: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hde3: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; // 
            12'hde4: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hde5: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hde6: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hde7: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hde8: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hde9: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdea: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdeb: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdec: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hded: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdee: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdef: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdf0: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'hdf1: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //

            //default : char_line_pixels <= '0;
            
/*
            //code x38
            12'he00: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he01: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he02: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he03: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he04: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he05: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he06: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he07: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he08: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he09: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he0a: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he0b: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he0c: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he0d: char_line_pixels <= 50'b00000000000000000001111111111000000000000000000000; //
            12'he0e: char_line_pixels <= 50'b00000000000000000001111111111000000000000000000000; //
            12'he0f: char_line_pixels <= 50'b00000000000000000111110000111110000000000000000000; //
            12'he10: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'he11: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'he12: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'he13: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'he14: char_line_pixels <= 50'b00000000000000000111110000111110000000000000000000; //
            12'he15: char_line_pixels <= 50'b00000000000000000001111111111000000000000000000000; //
            12'he16: char_line_pixels <= 50'b00000000000000000001111111111000000000000000000000; //
            12'he17: char_line_pixels <= 50'b00000000000000000111110000111110000000000000000000; //
            12'he18: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'he19: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'he1a: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'he1b: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'he1c: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'he1d: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'he1e: char_line_pixels <= 50'b00000000000000000111110000111110000000000000000000; //
            12'he1f: char_line_pixels <= 50'b00000000000000000001111111111000000000000000000000; //
            12'he20: char_line_pixels <= 50'b00000000000000000001111111111000000000000000000000; //
            12'he21: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he22: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he23: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; // 
            12'he24: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he25: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he26: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he27: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he28: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he29: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he2a: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he2b: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he2c: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he2d: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he2e: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he2f: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he30: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he31: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //


            //code x39
            12'he40: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he41: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he42: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he43: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he44: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he45: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he46: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he47: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he48: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he49: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he4a: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he4b: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he4c: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he4d: char_line_pixels <= 50'b00000000000000000001111111111000000000000000000000; //
            12'he4e: char_line_pixels <= 50'b00000000000000000001111111111000000000000000000000; //
            12'he4f: char_line_pixels <= 50'b00000000000000000111110000111110000000000000000000; //
            12'he50: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'he51: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'he52: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'he53: char_line_pixels <= 50'b00000000000000000111100000011110000000000000000000; //
            12'he54: char_line_pixels <= 50'b00000000000000000111110000111110000000000000000000; //
            12'he55: char_line_pixels <= 50'b00000000000000000011111111111110000000000000000000; //
            12'he56: char_line_pixels <= 50'b00000000000000000000111111111110000000000000000000; //
            12'he57: char_line_pixels <= 50'b00000000000000000000000000111110000000000000000000; //
            12'he58: char_line_pixels <= 50'b00000000000000000000000000011110000000000000000000; //
            12'he59: char_line_pixels <= 50'b00000000000000000000000000011110000000000000000000; //
            12'he5a: char_line_pixels <= 50'b00000000000000000000000000011110000000000000000000; //
            12'he5b: char_line_pixels <= 50'b00000000000000000000000000011110000000000000000000; //
            12'he5c: char_line_pixels <= 50'b00000000000000000000000000011110000000000000000000; //
            12'he5d: char_line_pixels <= 50'b00000000000000000000000000011110000000000000000000; //
            12'he5e: char_line_pixels <= 50'b00000000000000000000000000111110000000000000000000; //
            12'he5f: char_line_pixels <= 50'b00000000000000000001111111111000000000000000000000; //
            12'he60: char_line_pixels <= 50'b00000000000000000001111111111000000000000000000000; //
            12'he61: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he62: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he63: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; // 
            12'he64: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he65: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he66: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he67: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he68: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he69: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he6a: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he6b: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he6c: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he6d: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he6e: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he6f: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he70: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            12'he71: char_line_pixels <= 50'b00000000000000000000000000000000000000000000000000; //
            */
            
        endcase
    end

endmodule
