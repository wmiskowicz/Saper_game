`timescale 1ns / 1ps
// ROM with synchonous read (inferring Block RAM)
// character ROM
//  - 8-by-16 (8-by-2^4) font
//  - 128 (2^7) characters
//  - ROM size: 512-by-8 (2^11-by-8) bits
//              16K bits: 1 BRAM

module num_font_rom
    (
        input  wire        clk,
        input  wire [12:0] addr,            // {char_code[6:0], char_line[5:0]}
        output reg  [49:0]  char_line_pixels // pixels of the character line
    );

    // signal declaration
    reg [49:0] data;

    // body
    always @(posedge clk)
        char_line_pixels <= data;

    always @*
        case (addr)
            //code x00
            13'h000: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h001: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h002: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h003: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h004: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h005: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h006: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h007: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h008: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h009: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h00a: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h00b: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h00c: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h00d: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h00e: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h00f: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h010: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h011: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h012: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h013: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h014: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h015: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h016: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h017: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h018: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h019: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h01a: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h01b: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h01c: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h01d: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h01e: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h01f: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h020: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h021: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h022: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h023: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h024: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h025: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h026: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h027: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h028: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h029: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h02a: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h02b: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h02c: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h02d: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h02e: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h02f: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h030: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h031: data = 50'b00000000000000000000000000000000000000000000000000; //
            
            //code x03
            13'h0c0: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0c1: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0c2: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0c3: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0c4: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0c5: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0c6: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0c7: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0c8: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0c9: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0ca: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0cb: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0cc: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0cd: data = 50'b00000000000000000001110000111000000000000000000000;
            13'h0ce: data = 50'b00000000000000000011111001111100000000000000000000; //
            13'h0cf: data = 50'b00000000000000000111111111111110000000000000000000; //
            13'h0d0: data = 50'b00000000000000000111111111111110000000000000000000; //
            13'h0d1: data = 50'b00000000000000000111111111111110000000000000000000; //
            13'h0d2: data = 50'b00000000000000000111111111111110000000000000000000; //
            13'h0d3: data = 50'b00000000000000000111111111111110000000000000000000; //
            13'h0d4: data = 50'b00000000000000000111111111111110000000000000000000; //
            13'h0d5: data = 50'b00000000000000000111111111111110000000000000000000; //
            13'h0d6: data = 50'b00000000000000000111111111111110000000000000000000; //
            13'h0d7: data = 50'b00000000000000000011111111111100000000000000000000; //
            13'h0d8: data = 50'b00000000000000000001111111111000000000000000000000; //
            13'h0d9: data = 50'b00000000000000000000111111110000000000000000000000; //
            13'h0da: data = 50'b00000000000000000000011111100000000000000000000000; //
            13'h0db: data = 50'b00000000000000000000001111000000000000000000000000; //
            13'h0dc: data = 50'b00000000000000000000000110000000000000000000000000; //
            13'h0dd: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0de: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0df: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0e0: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0e1: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0e2: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0e3: data = 50'b00000000000000000000000000000000000000000000000000; // 
            13'h0e4: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0e5: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0e6: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0e7: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0e8: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0e9: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0ea: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0eb: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0ec: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0ed: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0ee: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0ef: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0f0: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'h0f1: data = 50'b00000000000000000000000000000000000000000000000000; //
  
            //code x30
            13'hc00: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc01: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc02: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc03: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc04: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc05: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc06: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc07: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc08: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc09: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc0a: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc0b: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc0c: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc0d: data = 50'b00000000000000000001111111111000000000000000000000;
            13'hc0e: data = 50'b00000000000000000001111111111000000000000000000000; //
            13'hc0f: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'hc10: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'hc11: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'hc12: data = 50'b00000000000000000111100000111110000000000000000000; //
            13'hc13: data = 50'b00000000000000000111100001111110000000000000000000; //
            13'hc14: data = 50'b00000000000000000111100011111110000000000000000000; //
            13'hc15: data = 50'b00000000000000000111100111111110000000000000000000; //
            13'hc16: data = 50'b00000000000000000111101111111110000000000000000000; //
            13'hc17: data = 50'b00000000000000000111111100011110000000000000000000; //
            13'hc18: data = 50'b00000000000000000111111000011110000000000000000000; //
            13'hc19: data = 50'b00000000000000000111110000011110000000000000000000; //
            13'hc1a: data = 50'b00000000000000000111110000011110000000000000000000; //
            13'hc1b: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'hc1c: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'hc1d: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'hc1e: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'hc1f: data = 50'b00000000000000000001111111111000000000000000000000; //
            13'hc20: data = 50'b00000000000000000001111111111000000000000000000000; //
            13'hc21: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc22: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc23: data = 50'b00000000000000000000000000000000000000000000000000; // 
            13'hc24: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc25: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc26: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc27: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc28: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc29: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc2a: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc2b: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc2c: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc2d: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc2e: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc2f: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc30: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc31: data = 50'b00000000000000000000000000000000000000000000000000; //


            //code x31
            13'hc40: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc41: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc42: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc43: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc44: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc45: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc46: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc47: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc48: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc49: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc4a: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc4b: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc4c: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc4d: data = 50'b00000000000000000000000111100000000000000000000000; //
            13'hc4e: data = 50'b00000000000000000000000111100000000000000000000000; //
            13'hc4f: data = 50'b00000000000000000000011111100000000000000000000000; //
            13'hc50: data = 50'b00000000000000000000011111100000000000000000000000; //
            13'hc51: data = 50'b00000000000000000001111111100000000000000000000000; //
            13'hc52: data = 50'b00000000000000000001111111100000000000000000000000; //
            13'hc53: data = 50'b00000000000000000000000111100000000000000000000000; //
            13'hc54: data = 50'b00000000000000000000000111100000000000000000000000; //
            13'hc55: data = 50'b00000000000000000000000111100000000000000000000000; //
            13'hc56: data = 50'b00000000000000000000000111100000000000000000000000; //
            13'hc57: data = 50'b00000000000000000000000111100000000000000000000000; //
            13'hc58: data = 50'b00000000000000000000000111100000000000000000000000; //
            13'hc59: data = 50'b00000000000000000000000111100000000000000000000000; //
            13'hc5a: data = 50'b00000000000000000000000111100000000000000000000000; //
            13'hc5b: data = 50'b00000000000000000000000111100000000000000000000000; //
            13'hc5c: data = 50'b00000000000000000000000111100000000000000000000000; //
            13'hc5d: data = 50'b00000000000000000000000111100000000000000000000000; //
            13'hc5e: data = 50'b00000000000000000000000111100000000000000000000000; //
            13'hc5f: data = 50'b00000000000000000000111111111100000000000000000000; //
            13'hc60: data = 50'b00000000000000000001111111111110000000000000000000; //
            13'hc61: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc62: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc63: data = 50'b00000000000000000000000000000000000000000000000000; // 
            13'hc64: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc65: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc66: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc67: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc68: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc69: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc6a: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc6b: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc6c: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc6d: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc6e: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc6f: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc70: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc71: data = 50'b00000000000000000000000000000000000000000000000000; //


            //code x32
            13'hc80: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc81: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc82: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc83: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc84: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc85: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc86: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc87: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc88: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc89: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc8a: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc8b: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc8c: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc8d: data = 50'b00000000000000000001111111111000000000000000000000; //
            13'hc8e: data = 50'b00000000000000000011111111111100000000000000000000; //
            13'hc8f: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'hc90: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'hc91: data = 50'b00000000000000000000000000011110000000000000000000; //
            13'hc92: data = 50'b00000000000000000000000000111100000000000000000000; //
            13'hc93: data = 50'b00000000000000000000000001111000000000000000000000; //
            13'hc94: data = 50'b00000000000000000000000011110000000000000000000000; //
            13'hc95: data = 50'b00000000000000000000000111100000000000000000000000; //
            13'hc96: data = 50'b00000000000000000000001111000000000000000000000000; //
            13'hc97: data = 50'b00000000000000000000011110000000000000000000000000; //
            13'hc98: data = 50'b00000000000000000000111100000000000000000000000000; //
            13'hc99: data = 50'b00000000000000000001111000000000000000000000000000; //
            13'hc9a: data = 50'b00000000000000000011110000000000000000000000000000; //
            13'hc9b: data = 50'b00000000000000000111100000000000000000000000000000; //
            13'hc9c: data = 50'b00000000000000000111100000000000000000000000000000; //
            13'hc9d: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'hc9e: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'hc9f: data = 50'b00000000000000000111111111111110000000000000000000; //
            13'hca0: data = 50'b00000000000000000111111111111110000000000000000000; //
            13'hca1: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hca2: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hca3: data = 50'b00000000000000000000000000000000000000000000000000; // 
            13'hca4: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hca5: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hca6: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hca7: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hca8: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hca9: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hcaa: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hcab: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hcac: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hcad: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hcae: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hcaf: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hcb0: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hcb1: data = 50'b00000000000000000000000000000000000000000000000000; //


            //code x33
            13'hc00: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc01: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc02: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc03: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc04: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc05: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc06: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc07: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc08: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc09: data = 50'b11000000000000000000000000000000000000000000000000; //
            13'hc0a: data = 50'b11000000000000000000000000000000000000000000000000; //
            13'hc0b: data = 50'b11000000000000000000000000000000000000000000000000; //
            13'hc0c: data = 50'b11000000000000000000000000000000000000000000000000; //
            13'hc0d: data = 50'b11000000000000000001111111111000000000000000000000; //
            13'hc0e: data = 50'b11000000000000000011111111111100000000000000000000; //
            13'hc0f: data = 50'b11000000000000000111100000011110000000000000000000; //
            13'hc10: data = 50'b11000000000000000111100000011110000000000000000000; //
            13'hc11: data = 50'b11000000000000000000000000011110000000000000000000; //
            13'hc12: data = 50'b11000000000000000000000000011110000000000000000000; //
            13'hc13: data = 50'b11000000000000000000000000011110000000000000000000; //
            13'hc14: data = 50'b11000000000000000000000000111100000000000000000000; //
            13'hc15: data = 50'b11000000000000000000011111111000000000000000000000; //
            13'hc16: data = 50'b11000000000000000000011111111000000000000000000000; //
            13'hc17: data = 50'b11000000000000000000000000111100000000000000000000; //
            13'hc18: data = 50'b11000000000000000000000000011110000000000000000000; //
            13'hc19: data = 50'b11000000000000000000000000011110000000000000000000; //
            13'hc1a: data = 50'b11000000000000000000000000011110000000000000000000; //
            13'hc1b: data = 50'b11000000000000000000000000011110000000000000000000; //
            13'hc1c: data = 50'b11000000000000000000000000011110000000000000000000; //
            13'hc1d: data = 50'b11000000000000000111100000011110000000000000000000; //
            13'hc1e: data = 50'b11000000000000000111100000011110000000000000000000; //
            13'hc1f: data = 50'b11000000000000000011111111111100000000000000000000; //
            13'hc20: data = 50'b11000000000000000001111111111000000000000000000000; //
            13'hc21: data = 50'b11000000000000000000000000000000000000000000000000; //
            13'hc22: data = 50'b11000000000000000000000000000000000000000000000000; //
            13'hc23: data = 50'b11000000000000000000000000000000000000000000000000; // 
            13'hc24: data = 50'b11000000000000000000000000000000000000000000000000; //
            13'hc25: data = 50'b11000000000000000000000000000000000000000000000000; //
            13'hc26: data = 50'b11000000000000000000000000000000000000000000000000; //
            13'hc27: data = 50'b11000000000000000000000000000000000000000000000000; //
            13'hc28: data = 50'b11000000000000000000000000000000000000000000000000; //
            13'hc29: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc2a: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc2b: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc2c: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc2d: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc2e: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc2f: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc30: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hc31: data = 50'b00000000000000000000000000000000000000000000000000; //


            //code x34
            13'hd00: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd01: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd02: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd03: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd04: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd05: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd06: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd07: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd08: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd09: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd0a: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd0b: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd0c: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd0d: data = 50'b00000000000000000000000000111000000000000000000000; //
            13'hd0e: data = 50'b00000000000000000000000001111000000000000000000000; //
            13'hd0f: data = 50'b00000000000000000000000111111000000000000000000000; //
            13'hd10: data = 50'b00000000000000000000000111111000000000000000000000; //
            13'hd11: data = 50'b00000000000000000000011111111000000000000000000000; //
            13'hd12: data = 50'b00000000000000000000011111111000000000000000000000; //
            13'hd13: data = 50'b00000000000000000001111001111000000000000000000000; //
            13'hd14: data = 50'b00000000000000000001111001111000000000000000000000; //
            13'hd15: data = 50'b00000000000000000111100001111000000000000000000000; //
            13'hd16: data = 50'b00000000000000000111100001111000000000000000000000; //
            13'hd17: data = 50'b00000000000000000111111111111110000000000000000000; //
            13'hd18: data = 50'b00000000000000000111111111111110000000000000000000; //
            13'hd19: data = 50'b00000000000000000000000001111000000000000000000000; //
            13'hd1a: data = 50'b00000000000000000000000001111000000000000000000000; //
            13'hd1b: data = 50'b00000000000000000000000001111000000000000000000000; //
            13'hd1c: data = 50'b00000000000000000000000001111000000000000000000000; //
            13'hd1d: data = 50'b00000000000000000000000001111000000000000000000000; //
            13'hd1e: data = 50'b00000000000000000000000001111000000000000000000000; //
            13'hd1f: data = 50'b00000000000000000000000011111100000000000000000000; //
            13'hd20: data = 50'b00000000000000000000000111111110000000000000000000; //
            13'hd21: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd22: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd23: data = 50'b00000000000000000000000000000000000000000000000000; // 
            13'hd24: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd25: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd26: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd27: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd28: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd29: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd2a: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd2b: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd2c: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd2d: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd2e: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd2f: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd30: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd31: data = 50'b00000000000000000000000000000000000000000000000000; //


            //code x35
            13'hd40: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd41: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd42: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd43: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd44: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd45: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd46: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd47: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd48: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd49: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd4a: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd4b: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd4c: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd4d: data = 50'b00000000000000000111111111111110000000000000000000; //
            13'hd4e: data = 50'b00000000000000000111111111111110000000000000000000; //
            13'hd4f: data = 50'b00000000000000000111100000000000000000000000000000; //
            13'hd50: data = 50'b00000000000000000111100000000000000000000000000000; //
            13'hd51: data = 50'b00000000000000000111100000000000000000000000000000; //
            13'hd52: data = 50'b00000000000000000111100000000000000000000000000000; //
            13'hd53: data = 50'b00000000000000000111100000000000000000000000000000; //
            13'hd54: data = 50'b00000000000000000111100000000000000000000000000000; //
            13'hd55: data = 50'b00000000000000000111111111110000000000000000000000; //
            13'hd56: data = 50'b00000000000000000011111111111100000000000000000000; //
            13'hd57: data = 50'b00000000000000000000000000011110000000000000000000; //
            13'hd58: data = 50'b00000000000000000000000000011110000000000000000000; //
            13'hd59: data = 50'b00000000000000000000000000011110000000000000000000; //
            13'hd5a: data = 50'b00000000000000000000000000011110000000000000000000; //
            13'hd5b: data = 50'b00000000000000000000000000011110000000000000000000; //
            13'hd5c: data = 50'b00000000000000000000000000011110000000000000000000; //
            13'hd5d: data = 50'b00000000000000000111000000011110000000000000000000; //
            13'hd5e: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'hd5f: data = 50'b00000000000000000011111111111000000000000000000000; //
            13'hd60: data = 50'b00000000000000000001111111110000000000000000000000; //
            13'hd61: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd62: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd63: data = 50'b00000000000000000000000000000000000000000000000000; // 
            13'hd64: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd65: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd66: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd67: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd68: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd69: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd6a: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd6b: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd6c: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd6d: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd6e: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd6f: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd70: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd71: data = 50'b00000000000000000000000000000000000000000000000000; //


            //code x36
            13'hd40: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd41: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd42: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd43: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd44: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd45: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd46: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd47: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd48: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd49: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd4a: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd4b: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd4c: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd4d: data = 50'b00000000000000000000001111110000000000000000000000; //
            13'hd4e: data = 50'b00000000000000000000111111100000000000000000000000; //
            13'hd4f: data = 50'b00000000000000000001111100000000000000000000000000; //
            13'hd50: data = 50'b00000000000000000011111000000000000000000000000000; //
            13'hd51: data = 50'b00000000000000000111110000000000000000000000000000; //
            13'hd52: data = 50'b00000000000000000111100000000000000000000000000000; //
            13'hd53: data = 50'b00000000000000000111100000000000000000000000000000; //
            13'hd54: data = 50'b00000000000000000111100000000000000000000000000000; //
            13'hd55: data = 50'b00000000000000000111111111111000000000000000000000; //
            13'hd56: data = 50'b00000000000000000111111111111100000000000000000000; //
            13'hd57: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'hd58: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'hd59: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'hd5a: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'hd5b: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'hd5c: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'hd5d: data = 50'b00000000000000000111000000011110000000000000000000; //
            13'hd5e: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'hd5f: data = 50'b00000000000000000011111111111100000000000000000000; //
            13'hd60: data = 50'b00000000000000000001111111110000000000000000000000; //
            13'hd61: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd62: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd63: data = 50'b00000000000000000000000000000000000000000000000000; // 
            13'hd64: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd65: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd66: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd67: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd68: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd69: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd6a: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd6b: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd6c: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd6d: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd6e: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd6f: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd70: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hd71: data = 50'b00000000000000000000000000000000000000000000000000; //


            //code x37
            13'hdc0: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hdc1: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hdc2: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hdc3: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hdc4: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hdc5: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hdc6: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hdc7: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hdc8: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hdc9: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hdca: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hdcb: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hdcc: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hdcd: data = 50'b00000000000000000111111111111110000000000000000000; //
            13'hdce: data = 50'b00000000000000000111111111111110000000000000000000; //
            13'hdcf: data = 50'b00000000000000000111110000111110000000000000000000; //
            13'hdd0: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'hdd1: data = 50'b00000000000000000000000000011110000000000000000000; //
            13'hdd2: data = 50'b00000000000000000000000000011110000000000000000000; //
            13'hdd3: data = 50'b00000000000000000000000000011110000000000000000000; //
            13'hdd4: data = 50'b00000000000000000000000000011110000000000000000000; //
            13'hdd5: data = 50'b000000000000000000000000000111100000000000000000000; //
            13'hdd6: data = 50'b00000000000000000000000001111000000000000000000000; //
            13'hdd7: data = 50'b00000000000000000000000111100000000000000000000000; //
            13'hdd8: data = 50'b00000000000000000000001111000000000000000000000000; //
            13'hdd9: data = 50'b00000000000000000000011110000000000000000000000000; //
            13'hdda: data = 50'b00000000000000000000011110000000000000000000000000; //
            13'hddb: data = 50'b00000000000000000000011110000000000000000000000000; //
            13'hddc: data = 50'b00000000000000000000011110000000000000000000000000; //
            13'hddd: data = 50'b00000000000000000000011110000000000000000000000000; //
            13'hdde: data = 50'b00000000000000000000011110000000000000000000000000; //
            13'hddf: data = 50'b00000000000000000000011110000000000000000000000000; //
            13'hde0: data = 50'b00000000000000000000011110000000000000000000000000; //
            13'hde1: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hde2: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hde3: data = 50'b00000000000000000000000000000000000000000000000000; // 
            13'hde4: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hde5: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hde6: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hde7: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hde8: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hde9: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hdea: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hdeb: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hdec: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hded: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hdee: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hdef: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hdf0: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'hdf1: data = 50'b00000000000000000000000000000000000000000000000000; //


            //code x38
            13'he00: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he01: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he02: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he03: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he04: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he05: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he06: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he07: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he08: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he09: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he0a: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he0b: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he0c: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he0d: data = 50'b00000000000000000001111111111000000000000000000000; //
            13'he0e: data = 50'b00000000000000000001111111111000000000000000000000; //
            13'he0f: data = 50'b00000000000000000111110000111110000000000000000000; //
            13'he10: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'he11: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'he12: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'he13: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'he14: data = 50'b00000000000000000111110000111110000000000000000000; //
            13'he15: data = 50'b00000000000000000001111111111000000000000000000000; //
            13'he16: data = 50'b00000000000000000001111111111000000000000000000000; //
            13'he17: data = 50'b00000000000000000111110000111110000000000000000000; //
            13'he18: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'he19: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'he1a: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'he1b: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'he1c: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'he1d: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'he1e: data = 50'b00000000000000000111110000111110000000000000000000; //
            13'he1f: data = 50'b00000000000000000001111111111000000000000000000000; //
            13'he20: data = 50'b00000000000000000001111111111000000000000000000000; //
            13'he21: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he22: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he23: data = 50'b00000000000000000000000000000000000000000000000000; // 
            13'he24: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he25: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he26: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he27: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he28: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he29: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he2a: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he2b: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he2c: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he2d: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he2e: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he2f: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he30: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he31: data = 50'b00000000000000000000000000000000000000000000000000; //


            //code x39
            13'he40: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he41: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he42: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he43: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he44: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he45: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he46: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he47: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he48: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he49: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he4a: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he4b: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he4c: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he4d: data = 50'b00000000000000000001111111111000000000000000000000; //
            13'he4e: data = 50'b00000000000000000001111111111000000000000000000000; //
            13'he4f: data = 50'b00000000000000000111110000111110000000000000000000; //
            13'he50: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'he51: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'he52: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'he53: data = 50'b00000000000000000111100000011110000000000000000000; //
            13'he54: data = 50'b00000000000000000111110000111110000000000000000000; //
            13'he55: data = 50'b00000000000000000011111111111110000000000000000000; //
            13'he56: data = 50'b00000000000000000000111111111110000000000000000000; //
            13'he57: data = 50'b00000000000000000000000000111110000000000000000000; //
            13'he58: data = 50'b00000000000000000000000000011110000000000000000000; //
            13'he59: data = 50'b00000000000000000000000000011110000000000000000000; //
            13'he5a: data = 50'b00000000000000000000000000011110000000000000000000; //
            13'he5b: data = 50'b00000000000000000000000000011110000000000000000000; //
            13'he5c: data = 50'b00000000000000000000000000011110000000000000000000; //
            13'he5d: data = 50'b00000000000000000000000000011110000000000000000000; //
            13'he5e: data = 50'b00000000000000000000000000111110000000000000000000; //
            13'he5f: data = 50'b00000000000000000001111111111000000000000000000000; //
            13'he60: data = 50'b00000000000000000001111111111000000000000000000000; //
            13'he61: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he62: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he63: data = 50'b00000000000000000000000000000000000000000000000000; // 
            13'he64: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he65: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he66: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he67: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he68: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he69: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he6a: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he6b: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he6c: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he6d: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he6e: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he6f: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he70: data = 50'b00000000000000000000000000000000000000000000000000; //
            13'he71: data = 50'b00000000000000000000000000000000000000000000000000; //
            
        endcase

endmodule
