`timescale 1ns / 1ps
// ROM with synchonous read (inferring Block RAM)
// character ROM
//  - 8-by-16 (8-by-2^4) font
//  - 128 (2^7) characters
//  - ROM size: 512-by-8 (2^11-by-8) bits
//              16K bits: 1 BRAM

module num_font_rom
    (
        input  wire        clk,
        input  wire [12:0] addr,            // {char_code[6:0], char_line[5:0]}
        output reg  [19:0]  char_line_pixels // pixels of the character line
    );

    // signal declaration
    reg [19:0] data;

    // body
    always @(posedge clk)
        char_line_pixels <= data;

    always @*
        case (addr)
            //code x00
            13'h000: data = 16'b00000000000000000000; //
            13'h001: data = 16'b00000000000000000000; //
            13'h002: data = 16'b00000000000000000000; //
            13'h003: data = 16'b00000000000000000000; //
            13'h004: data = 16'b00000000000000000000; //
            13'h005: data = 16'b00000000000000000000; //
            13'h006: data = 16'b00000000000000000000; //
            13'h007: data = 16'b00000000000000000000; //
            13'h008: data = 16'b00000000000000000000; //
            13'h009: data = 16'b00000000000000000000; //

            13'h00a: data = 16'b00000000000000000000; //
            13'h00b: data = 16'b00000000000000000000; //
            13'h00c: data = 16'b00000000000000000000; //
            13'h00d: data = 16'b00000000000000000000; //
            13'h00e: data = 16'b00000000000000000000; //
            13'h00f: data = 16'b00000000000000000000; //
            13'h010: data = 16'b00000000000000000000; //
            13'h011: data = 16'b00000000000000000000; //
            13'h012: data = 16'b00000000000000000000; //
            13'h013: data = 16'b00000000000000000000; //

            13'h014: data = 16'b00000000000000000000; //
            13'h015: data = 16'b00000000000000000000; //
            13'h016: data = 16'b00000000000000000000; //
            13'h017: data = 16'b00000000000000000000; //
            13'h018: data = 16'b00000000000000000000; //
            13'h019: data = 16'b00000000000000000000; //
            13'h01a: data = 16'b00000000000000000000; //
            13'h01b: data = 16'b00000000000000000000; //
            13'h01c: data = 16'b00000000000000000000; //
            13'h01d: data = 16'b00000000000000000000; //

            13'h01e: data = 16'b00000000000000000000; //
            13'h01f: data = 16'b00000000000000000000; //
            13'h020: data = 16'b00000000000000000000; //
            13'h021: data = 16'b00000000000000000000; //
            13'h022: data = 16'b00000000000000000000; //
            13'h023: data = 16'b00000000000000000000; //
            13'h024: data = 16'b00000000000000000000; //
            13'h025: data = 16'b00000000000000000000; //
            13'h026: data = 16'b00000000000000000000; //
            13'h027: data = 16'b00000000000000000000; //
            
            //code x03
            13'h030: data = 16'b00000000000000000000; //
            13'h031: data = 16'b00000000000000000000; //
            13'h032: data = 16'b00000000000000000000; //
            13'h033: data = 16'b00000000000000000000; //
            13'h034: data = 16'b01101100; //  ** **
            13'h035: data = 16'b11111110; // *******
            13'h036: data = 16'b11111110; // *******
            13'h037: data = 16'b11111110; // *******
            13'h038: data = 16'b11111110; // *******
            13'h039: data = 16'b01111100; //  *****
            13'h03a: data = 16'b00111000; //   ***
            13'h03b: data = 16'b00010000; //    *
            13'h03c: data = 16'b00000000000000000000; //
            13'h03d: data = 16'b00000000000000000000; //
            13'h03e: data = 16'b00000000000000000000; //
            13'h03f: data = 16'b00000000000000000000; //
            
           
          
  
            //code x30
            13'h300: data = 16'b00000000000000000000; //
            13'h301: data = 16'b00000000000000000000; //
            13'h302: data = 16'b01111100; //  *****
            13'h303: data = 16'b11000110; // **   **
            13'h304: data = 16'b11000110; // **   **
            13'h305: data = 16'b11001110; // **  ***
            13'h306: data = 16'b11011110; // ** ****
            13'h307: data = 16'b11110110; // **** **
            13'h308: data = 16'b11100110; // ***  **
            13'h309: data = 16'b11000110; // **   **
            13'h30a: data = 16'b11000110; // **   **
            13'h30b: data = 16'b01111100; //  *****
            13'h30c: data = 16'b00000000000000000000; //
            13'h30d: data = 16'b00000000000000000000; //
            13'h30e: data = 16'b00000000000000000000; //
            13'h30f: data = 16'b00000000000000000000; //
            //code x31
            13'h310: data = 16'b00000000000000000000; //
            13'h311: data = 16'b00000000000000000000; //
            13'h312: data = 16'b00011000; //
            13'h313: data = 16'b00111000; //
            13'h314: data = 16'b01111000; //    **
            13'h315: data = 16'b00011000; //   ***
            13'h316: data = 16'b00011000; //  ****
            13'h317: data = 16'b00011000; //    **
            13'h318: data = 16'b00011000; //    **
            13'h319: data = 16'b00011000; //    **
            13'h31a: data = 16'b00011000; //    **
            13'h31b: data = 16'b01111110; //    **
            13'h31c: data = 16'b00000000000000000000; //    **
            13'h31d: data = 16'b00000000000000000000; //  ******
            13'h31e: data = 16'b00000000000000000000; //
            13'h31f: data = 16'b00000000000000000000; //
            //code x32
            13'h320: data = 16'b00000000000000000000; //
            13'h321: data = 16'b00000000000000000000; //
            13'h322: data = 16'b01111100; //  *****
            13'h323: data = 16'b11000110; // **   **
            13'h324: data = 16'b00000110; //      **
            13'h325: data = 16'b00001100; //     **
            13'h326: data = 16'b00011000; //    **
            13'h327: data = 16'b00110000; //   **
            13'h328: data = 16'b01100000; //  **
            13'h329: data = 16'b11000000; // **
            13'h32a: data = 16'b11000110; // **   **
            13'h32b: data = 16'b11111110; // *******
            13'h32c: data = 16'b00000000000000000000; //
            13'h32d: data = 16'b00000000000000000000; //
            13'h32e: data = 16'b00000000000000000000; //
            13'h32f: data = 16'b00000000000000000000; //
            //code x33
            13'h330: data = 16'b00000000000000000000; //
            13'h331: data = 16'b00000000000000000000; //
            13'h332: data = 16'b01111100; //  *****
            13'h333: data = 16'b11000110; // **   **
            13'h334: data = 16'b00000110; //      **
            13'h335: data = 16'b00000110; //      **
            13'h336: data = 16'b00111100; //   ****
            13'h337: data = 16'b00000110; //      **
            13'h338: data = 16'b00000110; //      **
            13'h339: data = 16'b00000110; //      **
            13'h33a: data = 16'b11000110; // **   **
            13'h33b: data = 16'b01111100; //  *****
            13'h33c: data = 16'b00000000000000000000; //
            13'h33d: data = 16'b00000000000000000000; //
            13'h33e: data = 16'b00000000000000000000; //
            13'h33f: data = 16'b00000000000000000000; //
            //code x34
            13'h340: data = 16'b00000000000000000000; //
            13'h341: data = 16'b00000000000000000000; //
            13'h342: data = 16'b00001100; //     **
            13'h343: data = 16'b00011100; //    ***
            13'h344: data = 16'b00111100; //   ****
            13'h345: data = 16'b01101100; //  ** **
            13'h346: data = 16'b11001100; // **  **
            13'h347: data = 16'b11111110; // *******
            13'h348: data = 16'b00001100; //     **
            13'h349: data = 16'b00001100; //     **
            13'h34a: data = 16'b00001100; //     **
            13'h34b: data = 16'b00011110; //    ****
            13'h34c: data = 16'b00000000000000000000; //
            13'h34d: data = 16'b00000000000000000000; //
            13'h34e: data = 16'b00000000000000000000; //
            13'h34f: data = 16'b00000000000000000000; //
            //code x35
            13'h350: data = 16'b00000000000000000000; //
            13'h351: data = 16'b00000000000000000000; //
            13'h352: data = 16'b11111110; // *******
            13'h353: data = 16'b11000000; // **
            13'h354: data = 16'b11000000; // **
            13'h355: data = 16'b11000000; // **
            13'h356: data = 16'b11111100; // ******
            13'h357: data = 16'b00000110; //      **
            13'h358: data = 16'b00000110; //      **
            13'h359: data = 16'b00000110; //      **
            13'h35a: data = 16'b11000110; // **   **
            13'h35b: data = 16'b01111100; //  *****
            13'h35c: data = 16'b00000000000000000000; //
            13'h35d: data = 16'b00000000000000000000; //
            13'h35e: data = 16'b00000000000000000000; //
            13'h35f: data = 16'b00000000000000000000; //
            //code x36
            13'h360: data = 16'b00000000000000000000; //
            13'h361: data = 16'b00000000000000000000; //
            13'h362: data = 16'b00111000; //   ***
            13'h363: data = 16'b01100000; //  **
            13'h364: data = 16'b11000000; // **
            13'h365: data = 16'b11000000; // **
            13'h366: data = 16'b11111100; // ******
            13'h367: data = 16'b11000110; // **   **
            13'h368: data = 16'b11000110; // **   **
            13'h369: data = 16'b11000110; // **   **
            13'h36a: data = 16'b11000110; // **   **
            13'h36b: data = 16'b01111100; //  *****
            13'h36c: data = 16'b00000000000000000000; //
            13'h36d: data = 16'b00000000000000000000; //
            13'h36e: data = 16'b00000000000000000000; //
            13'h36f: data = 16'b00000000000000000000; //
            //code x37
            13'h370: data = 16'b00000000000000000000; //
            13'h371: data = 16'b00000000000000000000; //
            13'h372: data = 16'b11111110; // *******
            13'h373: data = 16'b11000110; // **   **
            13'h374: data = 16'b00000110; //      **
            13'h375: data = 16'b00000110; //      **
            13'h376: data = 16'b00001100; //     **
            13'h377: data = 16'b00011000; //    **
            13'h378: data = 16'b00110000; //   **
            13'h379: data = 16'b00110000; //   **
            13'h37a: data = 16'b00110000; //   **
            13'h37b: data = 16'b00110000; //   **
            13'h37c: data = 16'b00000000000000000000; //
            13'h37d: data = 16'b00000000000000000000; //
            13'h37e: data = 16'b00000000000000000000; //
            13'h37f: data = 16'b00000000000000000000; //
            //code x38
            13'h380: data = 16'b00000000000000000000; //
            13'h381: data = 16'b00000000000000000000; //
            13'h382: data = 16'b01111100; //  *****
            13'h383: data = 16'b11000110; // **   **
            13'h384: data = 16'b11000110; // **   **
            13'h385: data = 16'b11000110; // **   **
            13'h386: data = 16'b01111100; //  *****
            13'h387: data = 16'b11000110; // **   **
            13'h388: data = 16'b11000110; // **   **
            13'h389: data = 16'b11000110; // **   **
            13'h38a: data = 16'b11000110; // **   **
            13'h38b: data = 16'b01111100; //  *****
            13'h38c: data = 16'b00000000000000000000; //
            13'h38d: data = 16'b00000000000000000000; //
            13'h38e: data = 16'b00000000000000000000; //
            13'h38f: data = 16'b00000000000000000000; //
            //code x39
            13'h390: data = 16'b00000000000000000000; //
            13'h391: data = 16'b00000000000000000000; //
            13'h392: data = 16'b01111100; //  *****
            13'h393: data = 16'b11000110; // **   **
            13'h394: data = 16'b11000110; // **   **
            13'h395: data = 16'b11000110; // **   **
            13'h396: data = 16'b01111110; //  ******
            13'h397: data = 16'b00000110; //      **
            13'h398: data = 16'b00000110; //      **
            13'h399: data = 16'b00000110; //      **
            13'h39a: data = 16'b00001100; //     **
            13'h39b: data = 16'b01111000; //  ****
            13'h39c: data = 16'b00000000000000000000; //
            13'h39d: data = 16'b00000000000000000000; //
            13'h39e: data = 16'b00000000000000000000; //
            13'h39f: data = 16'b00000000000000000000; //
            
            
            
            
        endcase

endmodule
