/**
 * Copyright (C) 2023  AGH University of Science and Technology
 * MTM UEC2 Projekt
 * Author: Wojciech Miskowicz
 * 
 * Description:
 * Package with vga related constants.
 */

 package colour_pkg;

    // Parameters for drawing board, and button elements
    localparam [11:0] RED = 12'hf_0_0; 
    localparam [11:0] BLACK = 12'h1_1_1;
    
    localparam [11:0] BUTTON_BACK = 12'hd_d_d;
    localparam [11:0] BUTTON_WHITE = 12'hf_f_f;
    localparam [11:0] BUTTON_GRAY = 12'h5_5_5;
    
    endpackage
    