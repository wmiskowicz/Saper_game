`timescale 1ns / 1ps
// ROM with synchonous read (inferring Block RAM)
// character ROM
//  - 8-by-16 (8-by-2^4) font
//  - 128 (2^7) characters
//  - ROM size: 512-by-8 (2^11-by-8) bits
//              16K bits: 1 BRAM

module num_font_rom
    (
        input  wire        clk,
        input  wire [12:0] addr,            // {char_code[6:0], char_line[5:0]}
        output reg  [49:0]  char_line_pixels // pixels of the character line
    );

    // signal declaration
    reg [49:0] data;

    // body
    always @(posedge clk)
        char_line_pixels <= data;

    always @*
        case (addr)
            //code x00
            12'h000: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h001: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h002: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h003: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h004: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h005: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h006: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h007: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h008: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h009: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h00a: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h00b: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h00c: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h00d: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h00e: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h00f: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h010: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h011: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h012: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h013: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h014: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h015: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h016: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h017: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h018: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h019: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h01a: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h01b: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h01c: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h01d: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h01e: data = 50'b000000000000000000000000000000000000000000000000000000; //
            12'h01f: data = 50'b000000000000000000000000000000000000000000000000000000; //
            
            //code x03
            12'h060: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h061: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h062: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h063: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h064: data = 50'b00000000000000000001110000111000000000000000000000;
            12'h065: data = 50'b00000000000000000011111001111100000000000000000000; //
            12'h066: data = 50'b00000000000000000111111111111110000000000000000000; //
            12'h067: data = 50'b00000000000000000111111111111110000000000000000000; //
            12'h068: data = 50'b00000000000000000111111111111110000000000000000000; //
            12'h069: data = 50'b00000000000000000111111111111110000000000000000000; //
            12'h06a: data = 50'b00000000000000000111111111111110000000000000000000; //
            12'h06b: data = 50'b00000000000000000111111111111110000000000000000000; //
            12'h06c: data = 50'b00000000000000000111111111111110000000000000000000; //
            12'h06d: data = 50'b00000000000000000111111111111110000000000000000000; //
            12'h06e: data = 50'b00000000000000000011111111111100000000000000000000; //
            12'h06f: data = 50'b00000000000000000001111111111000000000000000000000; //
            12'h070: data = 50'b00000000000000000000111111110000000000000000000000; //
            12'h071: data = 50'b00000000000000000000011111100000000000000000000000; //
            12'h072: data = 50'b00000000000000000000001111000000000000000000000000; //
            12'h073: data = 50'b00000000000000000000000110000000000000000000000000; //
            12'h074: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h075: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h076: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h077: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h078: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h079: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h07a: data = 50'b00000000000000000000000000000000000000000000000000; // 
            12'h07b: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h07c: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h07d: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h07e: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h07f: data = 50'b00000000000000000000000000000000000000000000000000; //
  
            //code x30
            12'h600: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h601: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h602: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h603: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h604: data = 50'b00000000000000000001111111111000000000000000000000;
            12'h605: data = 50'b00000000000000000001111111111000000000000000000000; //
            12'h606: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h607: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h608: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h609: data = 50'b00000000000000000111100000111110000000000000000000; //
            12'h60a: data = 50'b00000000000000000111100001111110000000000000000000; //
            12'h60b: data = 50'b00000000000000000111100011111110000000000000000000; //
            12'h60c: data = 50'b00000000000000000111100111111110000000000000000000; //
            12'h60d: data = 50'b00000000000000000111101111111110000000000000000000; //
            12'h60e: data = 50'b00000000000000000111111100011110000000000000000000; //
            12'h60f: data = 50'b00000000000000000111111000011110000000000000000000; //
            12'h610: data = 50'b00000000000000000111110000011110000000000000000000; //
            12'h611: data = 50'b00000000000000000111110000011110000000000000000000; //
            12'h612: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h613: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h614: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h615: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h616: data = 50'b00000000000000000001111111111000000000000000000000; //
            12'h617: data = 50'b00000000000000000001111111111000000000000000000000; //
            12'h618: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h619: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h61a: data = 50'b00000000000000000000000000000000000000000000000000; // 
            12'h61b: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h61c: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h61d: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h61e: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h61f: data = 50'b00000000000000000000000000000000000000000000000000; //


            //code x31
            12'h620: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h621: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h622: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h623: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h624: data = 50'b00000000000000000000000111100000000000000000000000; //
            12'h625: data = 50'b00000000000000000000000111100000000000000000000000; //
            12'h626: data = 50'b00000000000000000000011111100000000000000000000000; //
            12'h627: data = 50'b00000000000000000000011111100000000000000000000000; //
            12'h628: data = 50'b00000000000000000001111111100000000000000000000000; //
            12'h629: data = 50'b00000000000000000001111111100000000000000000000000; //
            12'h62a: data = 50'b00000000000000000000000111100000000000000000000000; //
            12'h62b: data = 50'b00000000000000000000000111100000000000000000000000; //
            12'h62c: data = 50'b00000000000000000000000111100000000000000000000000; //
            12'h62d: data = 50'b00000000000000000000000111100000000000000000000000; //
            12'h62e: data = 50'b00000000000000000000000111100000000000000000000000; //
            12'h62f: data = 50'b00000000000000000000000111100000000000000000000000; //
            12'h630: data = 50'b00000000000000000000000111100000000000000000000000; //
            12'h631: data = 50'b00000000000000000000000111100000000000000000000000; //
            12'h632: data = 50'b00000000000000000000000111100000000000000000000000; //
            12'h633: data = 50'b00000000000000000000000111100000000000000000000000; //
            12'h634: data = 50'b00000000000000000000000111100000000000000000000000; //
            12'h635: data = 50'b00000000000000000000000111100000000000000000000000; //
            12'h636: data = 50'b00000000000000000000111111111100000000000000000000; //
            12'h637: data = 50'b00000000000000000001111111111110000000000000000000; //
            12'h638: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h639: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h63a: data = 50'b00000000000000000000000000000000000000000000000000; // 
            12'h63b: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h63c: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h63d: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h63e: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h63f: data = 50'b00000000000000000000000000000000000000000000000000; //


            //code x32
            12'h640: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h641: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h642: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h643: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h644: data = 50'b00000000000000000001111111111000000000000000000000; //
            12'h645: data = 50'b00000000000000000011111111111100000000000000000000; //
            12'h646: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h647: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h648: data = 50'b00000000000000000000000000011110000000000000000000; //
            12'h649: data = 50'b00000000000000000000000000111100000000000000000000; //
            12'h64a: data = 50'b00000000000000000000000001111000000000000000000000; //
            12'h64b: data = 50'b00000000000000000000000011110000000000000000000000; //
            12'h64c: data = 50'b00000000000000000000000111100000000000000000000000; //
            12'h64d: data = 50'b00000000000000000000001111000000000000000000000000; //
            12'h64e: data = 50'b00000000000000000000011110000000000000000000000000; //
            12'h64f: data = 50'b00000000000000000000111100000000000000000000000000; //
            12'h650: data = 50'b00000000000000000001111000000000000000000000000000; //
            12'h651: data = 50'b00000000000000000011110000000000000000000000000000; //
            12'h652: data = 50'b00000000000000000111100000000000000000000000000000; //
            12'h653: data = 50'b00000000000000000111100000000000000000000000000000; //
            12'h654: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h655: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h656: data = 50'b00000000000000000111111111111110000000000000000000; //
            12'h657: data = 50'b00000000000000000111111111111110000000000000000000; //
            12'h658: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h659: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h65a: data = 50'b00000000000000000000000000000000000000000000000000; // 
            12'h65b: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h65c: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h65d: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h65e: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h65f: data = 50'b00000000000000000000000000000000000000000000000000; //


            //code x33
            12'h660: data = 50'b11000000000000000000000000000000000000000000000000; //
            12'h661: data = 50'b11000000000000000000000000000000000000000000000000; //
            12'h662: data = 50'b11000000000000000000000000000000000000000000000000; //
            12'h663: data = 50'b11000000000000000000000000000000000000000000000000; //
            12'h664: data = 50'b11000000000000000001111111111000000000000000000000; //
            12'h665: data = 50'b11000000000000000011111111111100000000000000000000; //
            12'h666: data = 50'b11000000000000000111100000011110000000000000000000; //
            12'h667: data = 50'b11000000000000000111100000011110000000000000000000; //
            12'h668: data = 50'b11000000000000000000000000011110000000000000000000; //
            12'h669: data = 50'b11000000000000000000000000011110000000000000000000; //
            12'h66a: data = 50'b11000000000000000000000000011110000000000000000000; //
            12'h66b: data = 50'b11000000000000000000000000111100000000000000000000; //
            12'h66c: data = 50'b11000000000000000000011111111000000000000000000000; //
            12'h66d: data = 50'b11000000000000000000011111111000000000000000000000; //
            12'h66e: data = 50'b11000000000000000000000000111100000000000000000000; //
            12'h66f: data = 50'b11000000000000000000000000011110000000000000000000; //
            12'h670: data = 50'b11000000000000000000000000011110000000000000000000; //
            12'h671: data = 50'b11000000000000000000000000011110000000000000000000; //
            12'h672: data = 50'b11000000000000000000000000011110000000000000000000; //
            12'h673: data = 50'b11000000000000000000000000011110000000000000000000; //
            12'h674: data = 50'b11000000000000000111100000011110000000000000000000; //
            12'h675: data = 50'b11000000000000000111100000011110000000000000000000; //
            12'h676: data = 50'b11000000000000000011111111111100000000000000000000; //
            12'h677: data = 50'b11000000000000000001111111111000000000000000000000; //
            12'h678: data = 50'b11000000000000000000000000000000000000000000000000; //
            12'h679: data = 50'b11000000000000000000000000000000000000000000000000; //
            12'h67a: data = 50'b11000000000000000000000000000000000000000000000000; // 
            12'h67b: data = 50'b11000000000000000000000000000000000000000000000000; //
            12'h67c: data = 50'b11000000000000000000000000000000000000000000000000; //
            12'h67d: data = 50'b11000000000000000000000000000000000000000000000000; //
            12'h67e: data = 50'b11000000000000000000000000000000000000000000000000; //
            12'h67f: data = 50'b11000000000000000000000000000000000000000000000000; //


            //code x34
            12'h680: data = 50'b00000000000000000000000000000000000000000000000011; //
            12'h681: data = 50'b00000000000000000000000000000000000000000000000011; //
            12'h682: data = 50'b00000000000000000000000000000000000000000000000011; //
            12'h683: data = 50'b00000000000000000000000000000000000000000000000011; //
            12'h684: data = 50'b00000000000000000000000000111000000000000000000011; //
            12'h685: data = 50'b00000000000000000000000001111000000000000000000011; //
            12'h686: data = 50'b00000000000000000000000111111000000000000000000011; //
            12'h687: data = 50'b00000000000000000000000111111000000000000000000011; //
            12'h688: data = 50'b00000000000000000000011111111000000000000000000011; //
            12'h689: data = 50'b00000000000000000000011111111000000000000000000011; //
            12'h68a: data = 50'b00000000000000000001111001111000000000000000000011; //
            12'h68b: data = 50'b00000000000000000001111001111000000000000000000011; //
            12'h68c: data = 50'b00000000000000000111100001111000000000000000000011; //
            12'h68d: data = 50'b00000000000000000111100001111000000000000000000011; //
            12'h68e: data = 50'b00000000000000000111111111111110000000000000000011; //
            12'h68f: data = 50'b00000000000000000111111111111110000000000000000011; //
            12'h690: data = 50'b00000000000000000000000001111000000000000000000011; //
            12'h691: data = 50'b00000000000000000000000001111000000000000000000011; //
            12'h692: data = 50'b00000000000000000000000001111000000000000000000011; //
            12'h693: data = 50'b00000000000000000000000001111000000000000000000011; //
            12'h694: data = 50'b00000000000000000000000001111000000000000000000011; //
            12'h695: data = 50'b00000000000000000000000001111000000000000000000011; //
            12'h696: data = 50'b00000000000000000000000011111100000000000000000011; //
            12'h697: data = 50'b00000000000000000000000111111110000000000000000011; //
            12'h698: data = 50'b00000000000000000000000000000000000000000000000011; //
            12'h699: data = 50'b00000000000000000000000000000000000000000000000011; //
            12'h69a: data = 50'b00000000000000000000000000000000000000000000000011; // 
            12'h69b: data = 50'b00000000000000000000000000000000000000000000000011; //
            12'h69c: data = 50'b00000000000000000000000000000000000000000000000011; //
            12'h69d: data = 50'b00000000000000000000000000000000000000000000000011; //
            12'h69e: data = 50'b00000000000000000000000000000000000000000000000011; //
            12'h69f: data = 50'b00000000000000000000000000000000000000000000000011; //


            //code x35
            12'h6a0: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6a1: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6a2: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6a3: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6a4: data = 50'b00000000000000000111111111111110000000000000000000; //
            12'h6a5: data = 50'b00000000000000000111111111111110000000000000000000; //
            12'h6a6: data = 50'b00000000000000000111100000000000000000000000000000; //
            12'h6a7: data = 50'b00000000000000000111100000000000000000000000000000; //
            12'h6a8: data = 50'b00000000000000000111100000000000000000000000000000; //
            12'h6a9: data = 50'b00000000000000000111100000000000000000000000000000; //
            12'h6aa: data = 50'b00000000000000000111100000000000000000000000000000; //
            12'h6ab: data = 50'b00000000000000000111100000000000000000000000000000; //
            12'h6ac: data = 50'b00000000000000000111111111110000000000000000000000; //
            12'h6ad: data = 50'b00000000000000000011111111111100000000000000000000; //
            12'h6ae: data = 50'b00000000000000000000000000011110000000000000000000; //
            12'h6af: data = 50'b00000000000000000000000000011110000000000000000000; //
            12'h6b0: data = 50'b00000000000000000000000000011110000000000000000000; //
            12'h6b1: data = 50'b00000000000000000000000000011110000000000000000000; //
            12'h6b2: data = 50'b00000000000000000000000000011110000000000000000000; //
            12'h6b3: data = 50'b00000000000000000000000000011110000000000000000000; //
            12'h6b4: data = 50'b00000000000000000111000000011110000000000000000000; //
            12'h6b5: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h6b6: data = 50'b00000000000000000011111111111000000000000000000000; //
            12'h6b7: data = 50'b00000000000000000001111111110000000000000000000000; //
            12'h6b8: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6b9: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6ba: data = 50'b00000000000000000000000000000000000000000000000000; // 
            12'h6bb: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6bc: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6bd: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6be: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6bf: data = 50'b00000000000000000000000000000000000000000000000000; //


            //code x36
            12'h6c0: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6c1: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6c2: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6c3: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6c4: data = 50'b00000000000000000000001111110000000000000000000000; //
            12'h6c5: data = 50'b00000000000000000000111111100000000000000000000000; //
            12'h6c6: data = 50'b00000000000000000001111100000000000000000000000000; //
            12'h6c7: data = 50'b00000000000000000011111000000000000000000000000000; //
            12'h6c8: data = 50'b00000000000000000111110000000000000000000000000000; //
            12'h6c9: data = 50'b00000000000000000111100000000000000000000000000000; //
            12'h6ca: data = 50'b00000000000000000111100000000000000000000000000000; //
            12'h6cb: data = 50'b00000000000000000111100000000000000000000000000000; //
            12'h6cc: data = 50'b00000000000000000111111111111000000000000000000000; //
            12'h6cd: data = 50'b00000000000000000111111111111100000000000000000000; //
            12'h6ce: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h6cf: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h6d0: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h6d1: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h6d2: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h6d3: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h6d4: data = 50'b00000000000000000111000000011110000000000000000000; //
            12'h6d5: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h6d6: data = 50'b00000000000000000011111111111100000000000000000000; //
            12'h6d7: data = 50'b00000000000000000001111111110000000000000000000000; //
            12'h6d8: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6d9: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6da: data = 50'b00000000000000000000000000000000000000000000000000; // 
            12'h6db: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6dc: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6dd: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6de: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6df: data = 50'b00000000000000000000000000000000000000000000000000; //


            //code x37
            12'h6e0: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6e1: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6e2: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6e3: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6e4: data = 50'b00000000000000000111111111111110000000000000000000; //
            12'h6e5: data = 50'b00000000000000000111111111111110000000000000000000; //
            12'h6e6: data = 50'b00000000000000000111110000111110000000000000000000; //
            12'h6e7: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h6e8: data = 50'b00000000000000000000000000011110000000000000000000; //
            12'h6e9: data = 50'b00000000000000000000000000011110000000000000000000; //
            12'h6ea: data = 50'b00000000000000000000000000011110000000000000000000; //
            12'h6eb: data = 50'b00000000000000000000000000011110000000000000000000; //
            12'h6ec: data = 50'b000000000000000000000000000111100000000000000000000; //
            12'h6ed: data = 50'b00000000000000000000000001111000000000000000000000; //
            12'h6ee: data = 50'b00000000000000000000000111100000000000000000000000; //
            12'h6ef: data = 50'b00000000000000000000001111000000000000000000000000; //
            12'h6f0: data = 50'b00000000000000000000011110000000000000000000000000; //
            12'h6f1: data = 50'b00000000000000000000011110000000000000000000000000; //
            12'h6f2: data = 50'b00000000000000000000011110000000000000000000000000; //
            12'h6f3: data = 50'b00000000000000000000011110000000000000000000000000; //
            12'h6f4: data = 50'b00000000000000000000011110000000000000000000000000; //
            12'h6f5: data = 50'b00000000000000000000011110000000000000000000000000; //
            12'h6f6: data = 50'b00000000000000000000011110000000000000000000000000; //
            12'h6f7: data = 50'b00000000000000000000011110000000000000000000000000; //
            12'h6f8: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6f9: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6fa: data = 50'b00000000000000000000000000000000000000000000000000; // 
            12'h6fb: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6fc: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6fd: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6fe: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h6ff: data = 50'b00000000000000000000000000000000000000000000000000; //


            //code x38
            12'h700: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h701: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h702: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h703: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h704: data = 50'b00000000000000000001111111111000000000000000000000; //
            12'h705: data = 50'b00000000000000000001111111111000000000000000000000; //
            12'h706: data = 50'b00000000000000000111110000111110000000000000000000; //
            12'h707: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h708: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h709: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h70a: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h70b: data = 50'b00000000000000000111110000111110000000000000000000; //
            12'h70c: data = 50'b00000000000000000001111111111000000000000000000000; //
            12'h70d: data = 50'b00000000000000000001111111111000000000000000000000; //
            12'h70e: data = 50'b00000000000000000111110000111110000000000000000000; //
            12'h70f: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h710: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h711: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h712: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h713: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h714: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h715: data = 50'b00000000000000000111110000111110000000000000000000; //
            12'h716: data = 50'b00000000000000000001111111111000000000000000000000; //
            12'h717: data = 50'b00000000000000000001111111111000000000000000000000; //
            12'h718: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h719: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h71a: data = 50'b00000000000000000000000000000000000000000000000000; // 
            12'h71b: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h71c: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h71d: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h71e: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h71f: data = 50'b00000000000000000000000000000000000000000000000000; //


            //code x39
            12'h710: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h711: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h712: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h713: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h714: data = 50'b00000000000000000001111111111000000000000000000000; //
            12'h715: data = 50'b00000000000000000001111111111000000000000000000000; //
            12'h716: data = 50'b00000000000000000111110000111110000000000000000000; //
            12'h717: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h718: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h719: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h71a: data = 50'b00000000000000000111100000011110000000000000000000; //
            12'h71b: data = 50'b00000000000000000111110000111110000000000000000000; //
            12'h71c: data = 50'b00000000000000000011111111111110000000000000000000; //
            12'h71d: data = 50'b00000000000000000000111111111110000000000000000000; //
            12'h71e: data = 50'b00000000000000000000000000111110000000000000000000; //
            12'h71f: data = 50'b00000000000000000000000000011110000000000000000000; //
            12'h720: data = 50'b00000000000000000000000000011110000000000000000000; //
            12'h721: data = 50'b00000000000000000000000000011110000000000000000000; //
            12'h722: data = 50'b00000000000000000000000000011110000000000000000000; //
            12'h723: data = 50'b00000000000000000000000000011110000000000000000000; //
            12'h724: data = 50'b00000000000000000000000000011110000000000000000000; //
            12'h725: data = 50'b00000000000000000000000000111110000000000000000000; //
            12'h726: data = 50'b00000000000000000001111111111000000000000000000000; //
            12'h727: data = 50'b00000000000000000001111111111000000000000000000000; //
            12'h728: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h729: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h72a: data = 50'b00000000000000000000000000000000000000000000000000; // 
            12'h72b: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h72c: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h72d: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h72e: data = 50'b00000000000000000000000000000000000000000000000000; //
            12'h72f: data = 50'b00000000000000000000000000000000000000000000000000; //
            
        endcase

endmodule
