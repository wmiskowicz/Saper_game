`timescale 1ns / 1ps
// ROM with synchonous read (inferring Block RAM)
// character ROM
//  - 8-by-16 (8-by-2^4) font
//  - 128 (2^7) characters
//  - ROM size: 512-by-8 (2^11-by-8) bits
//              16K bits: 1 BRAM

module num_font_rom
    (
        input  wire        clk,
        input  wire [11:0] addr,            // {char_code[6:0], char_line[4:0]}
        output reg  [19:0]  char_line_pixels // pixels of the character line
    );

    // signal declaration
    reg [19:0] data;

    // body
    always @(posedge clk)
        char_line_pixels <= data;

    always @*
        case (addr)
            //code x00
            12'h000: data = 16'b00000000000000000000; //
            12'h001: data = 16'b00000000000000000000; //
            12'h002: data = 16'b00000000000000000000; //
            12'h003: data = 16'b00000000000000000000; //
            12'h004: data = 16'b00000000000000000000; //
            12'h005: data = 16'b00000000000000000000; //
            12'h006: data = 16'b00000000000000000000; //
            12'h007: data = 16'b00000000000000000000; //
            12'h008: data = 16'b00000000000000000000; //
            12'h009: data = 16'b00000000000000000000; //
            12'h00a: data = 16'b00000000000000000000; //
            12'h00b: data = 16'b00000000000000000000; //
            12'h00c: data = 16'b00000000000000000000; //
            12'h00d: data = 16'b00000000000000000000; //
            12'h00e: data = 16'b00000000000000000000; //
            12'h00f: data = 16'b00000000000000000000; //
            12'h010: data = 16'b00000000000000000000; //
            12'h011: data = 16'b00000000000000000000; //
            12'h012: data = 16'b00000000000000000000; //
            12'h013: data = 16'b00000000000000000000; //
            12'h014: data = 16'b00000000000000000000; //
            12'h015: data = 16'b00000000000000000000; //
            12'h016: data = 16'b00000000000000000000; //
            12'h017: data = 16'b00000000000000000000; //
            12'h018: data = 16'b00000000000000000000; //
            12'h019: data = 16'b00000000000000000000; //
            12'h01a: data = 16'b00000000000000000000; //
            12'h01b: data = 16'b00000000000000000000; //
            12'h01c: data = 16'b00000000000000000000; //
            12'h01d: data = 16'b00000000000000000000; //
            12'h01e: data = 16'b00000000000000000000; //
            12'h01f: data = 16'b00000000000000000000; //
            
            //code x03
            12'h000: data = 16'b0000000000000000; //
            12'h001: data = 16'b0000000000000000; //
            12'h002: data = 16'b0000000000000000; //
            12'h003: data = 16'b0000000000000000; //
            12'h004: data = 16'b0011100001110000;
            12'h005: data = 16'b0111110011111000; //
            12'h006: data = 16'b1111111111111100; //
            12'h007: data = 16'b1111111111111100; //
            12'h008: data = 16'b1111111111111100; //
            12'h009: data = 16'b1111111111111100; //
            12'h00a: data = 16'b1111111111111100; //
            12'h00b: data = 16'b1111111111111100; //
            12'h00c: data = 16'b1111111111111100; //
            12'h00d: data = 16'b1111111111111100; //
            12'h00e: data = 16'b0111111111111000; //
            12'h00f: data = 16'b0011111111110000; //
            12'h010: data = 16'b0001111111100000; //
            12'h011: data = 16'b0000111111000000; //
            12'h012: data = 16'b0000011110000000; //
            12'h013: data = 16'b0000001100000000; //
            12'h014: data = 16'b0000000000000000; //
            12'h015: data = 16'b0000000000000000; //
            12'h016: data = 16'b0000000000000000; //
            12'h017: data = 16'b0000000000000000; //
            12'h018: data = 16'b0000000000000000; //
            12'h019: data = 16'b0000000000000000; //
            12'h01a: data = 16'b0000000000000000; // 
            12'h01b: data = 16'b0000000000000000; //
            12'h01c: data = 16'b0000000000000000; //
            12'h01d: data = 16'b0000000000000000; //
            12'h01e: data = 16'b0000000000000000; //
            12'h01f: data = 16'b0000000000000000; //
  
            //code x30
            12'h000: data = 16'b0000000000000000; //
            12'h001: data = 16'b0000000000000000; //
            12'h002: data = 16'b0000000000000000; //
            12'h003: data = 16'b0000000000000000; //
            12'h004: data = 16'b0011111111110000;
            12'h005: data = 16'b0011111111110000; //
            12'h006: data = 16'b1111000000111100; //
            12'h007: data = 16'b1111000000111100; //
            12'h008: data = 16'b1111000000111100; //
            12'h009: data = 16'b1111000001111100; //
            12'h00a: data = 16'b1111000011111100; //
            12'h00b: data = 16'b1111000111111100; //
            12'h00c: data = 16'b1111001111111100; //
            12'h00d: data = 16'b1111011111111100; //
            12'h00e: data = 16'b1111111000111100; //
            12'h00f: data = 16'b1111110000111100; //
            12'h010: data = 16'b1111100000111100; //
            12'h011: data = 16'b1111100000111100; //
            12'h012: data = 16'b1111000000111100; //
            12'h013: data = 16'b1111000000111100; //
            12'h014: data = 16'b1111000000111100; //
            12'h015: data = 16'b1111000000111100; //
            12'h016: data = 16'b0011111111110000; //
            12'h017: data = 16'b0011111111110000; //
            12'h018: data = 16'b0000000000000000; //
            12'h019: data = 16'b0000000000000000; //
            12'h01a: data = 16'b0000000000000000; // 
            12'h01b: data = 16'b0000000000000000; //
            12'h01c: data = 16'b0000000000000000; //
            12'h01d: data = 16'b0000000000000000; //
            12'h01e: data = 16'b0000000000000000; //
            12'h01f: data = 16'b0000000000000000; //


            //code x31
            12'h000: data = 16'b0000000000000000; //
            12'h001: data = 16'b0000000000000000; //
            12'h002: data = 16'b0000000000000000; //
            12'h003: data = 16'b0000000000000000; //
            12'h004: data = 16'b0000001111000000; //
            12'h005: data = 16'b0000001111000000; //
            12'h006: data = 16'b0000111111000000; //
            12'h007: data = 16'b0000111111000000; //
            12'h008: data = 16'b0011111111000000; //
            12'h009: data = 16'b0011111111000000; //
            12'h00a: data = 16'b0000001111000000; //
            12'h00b: data = 16'b0000001111000000; //
            12'h00c: data = 16'b0000001111000000; //
            12'h00d: data = 16'b0000001111000000; //
            12'h00e: data = 16'b0000001111000000; //
            12'h00f: data = 16'b0000001111000000; //
            12'h010: data = 16'b0000001111000000; //
            12'h011: data = 16'b0000001111000000; //
            12'h012: data = 16'b0000001111000000; //
            12'h013: data = 16'b0000001111000000; //
            12'h014: data = 16'b0000001111000000; //
            12'h015: data = 16'b0000001111000000; //
            12'h016: data = 16'b0011111111111100; //
            12'h017: data = 16'b0011111111111100; //
            12'h018: data = 16'b0000000000000000; //
            12'h019: data = 16'b0000000000000000; //
            12'h01a: data = 16'b0000000000000000; // 
            12'h01b: data = 16'b0000000000000000; //
            12'h01c: data = 16'b0000000000000000; //
            12'h01d: data = 16'b0000000000000000; //
            12'h01e: data = 16'b0000000000000000; //
            12'h01f: data = 16'b0000000000000000; //


            //code x32
            12'h000: data = 16'b0000000000000000; //
            12'h001: data = 16'b0000000000000000; //
            12'h002: data = 16'b0000000000000000; //
            12'h003: data = 16'b0000000000000000; //
            12'h004: data = 16'b0011111111110000; //
            12'h005: data = 16'b0111111111111000; //
            12'h006: data = 16'b1111000000111100; //
            12'h007: data = 16'b1111000000111100; //
            12'h008: data = 16'b0000000000111100; //
            12'h009: data = 16'b0000000001111000; //
            12'h00a: data = 16'b0000000011110000; //
            12'h00b: data = 16'b0000000111100000; //
            12'h00c: data = 16'b0000001111000000; //
            12'h00d: data = 16'b0000011110000000; //
            12'h00e: data = 16'b0000111100000000; //
            12'h00f: data = 16'b0001111000000000; //
            12'h010: data = 16'b0011110000000000; //
            12'h011: data = 16'b0111100000000000; //
            12'h012: data = 16'b1111000000000000; //
            12'h013: data = 16'b1111000000000000; //
            12'h014: data = 16'b1111000000111100; //
            12'h015: data = 16'b1111000000111100; //
            12'h016: data = 16'b1111111111111100; //
            12'h017: data = 16'b1111111111111100; //
            12'h018: data = 16'b0000000000000000; //
            12'h019: data = 16'b0000000000000000; //
            12'h01a: data = 16'b0000000000000000; // 
            12'h01b: data = 16'b0000000000000000; //
            12'h01c: data = 16'b0000000000000000; //
            12'h01d: data = 16'b0000000000000000; //
            12'h01e: data = 16'b0000000000000000; //
            12'h01f: data = 16'b0000000000000000; //


            //code x33
            12'h000: data = 16'b0000000000000000; //
            12'h001: data = 16'b0000000000000000; //
            12'h002: data = 16'b0000000000000000; //
            12'h003: data = 16'b0000000000000000; //
            12'h004: data = 16'b0011111111110000; //
            12'h005: data = 16'b0111111111111000; //
            12'h006: data = 16'b1111000000111100; //
            12'h007: data = 16'b1111000000111100; //
            12'h008: data = 16'b0000000000111100; //
            12'h009: data = 16'b0000000000111100; //
            12'h00a: data = 16'b0000000000111100; //
            12'h00b: data = 16'b0000000001111000; //
            12'h00c: data = 16'00001111111110000; //
            12'h00d: data = 16'00001111111110000; //
            12'h00e: data = 16'b0000000001111000; //
            12'h00f: data = 16'b0000000000111100; //
            12'h010: data = 16'b0000000000111100; //
            12'h011: data = 16'b0000000000111100; //
            12'h012: data = 16'b0000000000111100; //
            12'h013: data = 16'b0000000000111100; //
            12'h014: data = 16'b1111000000111100; //
            12'h015: data = 16'b1111000000111100; //
            12'h016: data = 16'b0111111111111000; //
            12'h017: data = 16'b0011111111110000; //
            12'h018: data = 16'b0000000000000000; //
            12'h019: data = 16'b0000000000000000; //
            12'h01a: data = 16'b0000000000000000; // 
            12'h01b: data = 16'b0000000000000000; //
            12'h01c: data = 16'b0000000000000000; //
            12'h01d: data = 16'b0000000000000000; //
            12'h01e: data = 16'b0000000000000000; //
            12'h01f: data = 16'b0000000000000000; //


            //code x34
            12'h000: data = 16'b0000000000000000; //
            12'h001: data = 16'b0000000000000000; //
            12'h002: data = 16'b0000000000000000; //
            12'h003: data = 16'b0000000000000000; //
            12'h004: data = 16'b0000000001110000; //
            12'h005: data = 16'b0000000011110000; //
            12'h006: data = 16'b0000001111110000; //
            12'h007: data = 16'b0000001111110000; //
            12'h008: data = 16'b0000111111110000; //
            12'h009: data = 16'b0000111111110000; //
            12'h00a: data = 16'b0011110011110000; //
            12'h00b: data = 16'b0011110011110000; //
            12'h00c: data = 16'b1111000011110000; //
            12'h00d: data = 16'b1111000011110000; //
            12'h00e: data = 16'b1111111111111100; //
            12'h00f: data = 16'b1111111111111100; //
            12'h010: data = 16'b0000000011110000; //
            12'h011: data = 16'b0000000011110000; //
            12'h012: data = 16'b0000000011110000; //
            12'h013: data = 16'b0000000011110000; //
            12'h014: data = 16'b0000000011110000; //
            12'h015: data = 16'b0000000011110000; //
            12'h016: data = 16'b0000000111111000; //
            12'h017: data = 16'b0000001111111100; //
            12'h018: data = 16'b0000000000000000; //
            12'h019: data = 16'b0000000000000000; //
            12'h01a: data = 16'b0000000000000000; // 
            12'h01b: data = 16'b0000000000000000; //
            12'h01c: data = 16'b0000000000000000; //
            12'h01d: data = 16'b0000000000000000; //
            12'h01e: data = 16'b0000000000000000; //
            12'h01f: data = 16'b0000000000000000; //


            //code x35
            12'h000: data = 16'b0000000000000000; //
            12'h001: data = 16'b0000000000000000; //
            12'h002: data = 16'b0000000000000000; //
            12'h003: data = 16'b0000000000000000; //
            12'h004: data = 16'b1111111111111100; //
            12'h005: data = 16'b1111111111111100; //
            12'h006: data = 16'b1111000000000000; //
            12'h007: data = 16'b1111000000000000; //
            12'h008: data = 16'b1111000000000000; //
            12'h009: data = 16'b1111000000000000; //
            12'h00a: data = 16'b1111000000000000; //
            12'h00b: data = 16'b1111000000000000; //
            12'h00c: data = 16'b1111111111100000; //
            12'h00d: data = 16'b0111111111111000; //
            12'h00e: data = 16'b0000000000111100; //
            12'h00f: data = 16'b0000000000111100; //
            12'h010: data = 16'b0000000000111100; //
            12'h011: data = 16'b0000000000111100; //
            12'h012: data = 16'b0000000000111100; //
            12'h013: data = 16'b0000000000111100; //
            12'h014: data = 16'b1110000000111100; //
            12'h015: data = 16'b1111000000111100; //
            12'h016: data = 16'00111111111110000; //
            12'h017: data = 16'00011111111100000; //
            12'h018: data = 16'b0000000000000000; //
            12'h019: data = 16'b0000000000000000; //
            12'h01a: data = 16'b0000000000000000; // 
            12'h01b: data = 16'b0000000000000000; //
            12'h01c: data = 16'b0000000000000000; //
            12'h01d: data = 16'b0000000000000000; //
            12'h01e: data = 16'b0000000000000000; //
            12'h01f: data = 16'b0000000000000000; //


            //code x36
            12'h000: data = 16'b0000000000000000; //
            12'h001: data = 16'b0000000000000000; //
            12'h002: data = 16'b0000000000000000; //
            12'h003: data = 16'b0000000000000000; //
            12'h004: data = 16'b0000011111100000; //
            12'h005: data = 16'b0001111111000000; //
            12'h006: data = 16'b0011111000000000; //
            12'h007: data = 16'b0111110000000000; //
            12'h008: data = 16'b1111100000000000; //
            12'h009: data = 16'b1111000000000000; //
            12'h00a: data = 16'b1111000000000000; //
            12'h00b: data = 16'b1111000000000000; //
            12'h00c: data = 16'b1111111111110000; //
            12'h00d: data = 16'b1111111111111000; //
            12'h00e: data = 16'b1111000000111100; //
            12'h00f: data = 16'b1111000000111100; //
            12'h010: data = 16'b1111000000111100; //
            12'h011: data = 16'b1111000000111100; //
            12'h012: data = 16'b1111000000111100; //
            12'h013: data = 16'b1111000000111100; //
            12'h014: data = 16'b1110000000111100; //
            12'h015: data = 16'b1111000000111100; //
            12'h016: data = 16'00111111111111000; //
            12'h017: data = 16'00011111111100000; //
            12'h018: data = 16'b0000000000000000; //
            12'h019: data = 16'b0000000000000000; //
            12'h01a: data = 16'b0000000000000000; // 
            12'h01b: data = 16'b0000000000000000; //
            12'h01c: data = 16'b0000000000000000; //
            12'h01d: data = 16'b0000000000000000; //
            12'h01e: data = 16'b0000000000000000; //
            12'h01f: data = 16'b0000000000000000; //


            //code x37
            12'h000: data = 16'b0000000000000000; //
            12'h001: data = 16'b0000000000000000; //
            12'h002: data = 16'b0000000000000000; //
            12'h003: data = 16'b0000000000000000; //
            12'h004: data = 16'b1111111111111100; //
            12'h005: data = 16'b1111111111111100; //
            12'h006: data = 16'b1111100001111100; //
            12'h007: data = 16'b1111000000111100; //
            12'h008: data = 16'b0000000000111100; //
            12'h009: data = 16'b0000000000111100; //
            12'h00a: data = 16'b0000000000111100; //
            12'h00b: data = 16'b0000000000111100; //
            12'h00c: data = 16'b00000000001111000; //
            12'h00d: data = 16'b0000000011110000; //
            12'h00e: data = 16'b0000001111000000; //
            12'h00f: data = 16'b0000011110000000; //
            12'h010: data = 16'b0000111100000000; //
            12'h011: data = 16'b0000111100000000; //
            12'h012: data = 16'b0000111100000000; //
            12'h013: data = 16'b0000111100000000; //
            12'h014: data = 16'b0000111100000000; //
            12'h015: data = 16'b0000111100000000; //
            12'h016: data = 16'b0000111100000000; //
            12'h017: data = 16'b0000111100000000; //
            12'h018: data = 16'b0000000000000000; //
            12'h019: data = 16'b0000000000000000; //
            12'h01a: data = 16'b0000000000000000; // 
            12'h01b: data = 16'b0000000000000000; //
            12'h01c: data = 16'b0000000000000000; //
            12'h01d: data = 16'b0000000000000000; //
            12'h01e: data = 16'b0000000000000000; //
            12'h01f: data = 16'b0000000000000000; //


            //code x38
            12'h000: data = 16'b0000000000000000; //
            12'h001: data = 16'b0000000000000000; //
            12'h002: data = 16'b0000000000000000; //
            12'h003: data = 16'b0000000000000000; //
            12'h004: data = 16'b0011111111110000; //
            12'h005: data = 16'b0011111111110000; //
            12'h006: data = 16'b1111100001111100; //
            12'h007: data = 16'b1111000000111100; //
            12'h008: data = 16'b1111000000111100; //
            12'h009: data = 16'b1111000000111100; //
            12'h00a: data = 16'b1111000000111100; //
            12'h00b: data = 16'b1111100001111100; //
            12'h00c: data = 16'b0011111111110000; //
            12'h00d: data = 16'b0011111111110000; //
            12'h00e: data = 16'b1111100001111100; //
            12'h00f: data = 16'b1111000000111100; //
            12'h010: data = 16'b1111000000111100; //
            12'h011: data = 16'b1111000000111100; //
            12'h012: data = 16'b1111000000111100; //
            12'h013: data = 16'b1111000000111100; //
            12'h014: data = 16'b1111000000111100; //
            12'h015: data = 16'b1111100001111100; //
            12'h016: data = 16'b0011111111110000; //
            12'h017: data = 16'b0011111111110000; //
            12'h018: data = 16'b0000000000000000; //
            12'h019: data = 16'b0000000000000000; //
            12'h01a: data = 16'b0000000000000000; // 
            12'h01b: data = 16'b0000000000000000; //
            12'h01c: data = 16'b0000000000000000; //
            12'h01d: data = 16'b0000000000000000; //
            12'h01e: data = 16'b0000000000000000; //
            12'h01f: data = 16'b0000000000000000; //


            //code x39
            12'h000: data = 16'b0000000000000000; //
            12'h001: data = 16'b0000000000000000; //
            12'h002: data = 16'b0000000000000000; //
            12'h003: data = 16'b0000000000000000; //
            12'h004: data = 16'b0011111111110000; //
            12'h005: data = 16'b0011111111110000; //
            12'h006: data = 16'b1111100001111100; //
            12'h007: data = 16'b1111000000111100; //
            12'h008: data = 16'b1111000000111100; //
            12'h009: data = 16'b1111000000111100; //
            12'h00a: data = 16'b1111000000111100; //
            12'h00b: data = 16'b1111100001111100; //
            12'h00c: data = 16'b0111111111111100; //
            12'h00d: data = 16'b0001111111111100; //
            12'h00e: data = 16'b0000000001111100; //
            12'h00f: data = 16'b0000000000111100; //
            12'h010: data = 16'b0000000000111100; //
            12'h011: data = 16'b0000000000111100; //
            12'h012: data = 16'b0000000000111100; //
            12'h013: data = 16'b0000000000111100; //
            12'h014: data = 16'b0000000000111100; //
            12'h015: data = 16'b0000000001111100; //
            12'h016: data = 16'b0011111111110000; //
            12'h017: data = 16'b0011111111110000; //
            12'h018: data = 16'b0000000000000000; //
            12'h019: data = 16'b0000000000000000; //
            12'h01a: data = 16'b0000000000000000; // 
            12'h01b: data = 16'b0000000000000000; //
            12'h01c: data = 16'b0000000000000000; //
            12'h01d: data = 16'b0000000000000000; //
            12'h01e: data = 16'b0000000000000000; //
            12'h01f: data = 16'b0000000000000000; //
            
        endcase

endmodule
